

YPressurePump soln1 1 2 pressure=100k chemConcentration=100m
Ychannel soln1_channel 1 2 3 4 length=7.65m


Ychannel output0 5 0 6 7 length=5.9m
Ychannel connect1 8 9 10 11 length=1.18m
Ychannel connect2 12 13 14 15 length=1.18m
Ychannel connect3 16 17 18 19 length=2.15m
Ychannel connect4 20 21 22 23 length=3.27m
Ychannel connect5 24 25 26 27 length=15.05m
Yserpentine_50px_0 serp1 3 8 4 10
Yserpentine_150px_0 serp2 9 12 11 14
Yserpentine_300px_0 serp4 13 16 15 18
Yserpentine_300px_0 serp5 17 20 19 22
Yserpentine_300px_0 serp6 21 24 23 26
Yserpentine_300px_0 serp11 25 5 27 6


.tran 0.1m 1m
.print tran V(6)
.end


