

YPressurePump soln1 1 2 pressure=100k
Ychannel soln1_channel 1 3 2 4 length=7.65m

YPressurePump soln2 5 6 pressure=100k
Ychannel soln2_channel 5 7 6 8 length=3.24m

YPressurePump soln3 9 10 pressure=100k chemConcentration=100m
Ychannel soln3_channel 9 11 10 12 length=5.71m


Ychannel output0 13 0 14 15 length=5.9m
Ychannel connect1 16 17 18 19 length=1.18m
Ychannel connect2 20 21 22 23 length=1.18m
Ychannel connect3 24 25 26 27 length=2.15m
Ychannel connect4 28 29 30 31 length=3.27m
Ychannel connect5 32 33 34 35 length=15.05m
Ychannel connect6 36 37 38 39 length=4.41m
Ychannel connect7 40 41 42 43 length=2.68m
Yserpentine_50px_0 serp1 7 16 8 18
Yserpentine_150px_0 serp2 17 20 19 22
Ydiffmix_25px_0 mix0 3 21 24 4 23 26
Yserpentine_300px_0 serp3 11 28 12 30
Yserpentine_300px_0 serp4 29 32 31 34
Yserpentine_300px_0 serp5 33 36 35 38
Yserpentine_300px_0 serp6 37 44 39 45
Ydiffmix_25px_0 mix1 25 46 40 27 47 42
Yserpentine_300px_0 serp11 41 13 43 14


.tran 0.1m 1m


.end


